interface my_if(input clk, rstn);
  logic[7:0]data;
  logic valid;
endinterface
